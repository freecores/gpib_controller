--------------------------------------------------------------------------------
-- Entity: MemoryBlock
-- Date:2011-11-14  
-- Author: Administrator     
--
-- Description ${cursor}
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

library UNISIM;
use UNISIM.vcomponents.all;

use work.utilPkg.all;
use work.helperComponents.all;


entity MemoryBlock is
	port (
		reset : in std_logic;
		clk : in std_logic;
		-------------------------------------------------
		p1_addr : in std_logic_vector(10 downto 0);
		p1_data_in : in std_logic_vector(7 downto 0);
		p1_strobe : in std_logic;
		p1_data_out : out std_logic_vector(7 downto 0);
		-------------------------------------------------
		p2_addr : in std_logic_vector(10 downto 0);
		p2_data_in : in std_logic_vector(7 downto 0);
		p2_strobe : in std_logic;
		p2_data_out : out std_logic_vector(7 downto 0)
	);
end MemoryBlock;

architecture arch of MemoryBlock is

	constant ADDR_WIDTH : integer := 11;
	constant DATA_WIDTH : integer := 8;


	signal m_p1_parity_in, m_p1_parity_out : std_logic_vector(0 downto 0);
	signal m_p1_data_in, m_p1_data_out :
		std_logic_vector((DATA_WIDTH-1) downto 0);
	signal m_p1_addr : std_logic_vector((ADDR_WIDTH-1) downto 0);
	signal m_p1_clk, m_p1_en, m_p1_ssr, m_p1_we : std_logic;

	signal m_p2_parity_in, m_p2_parity_out : std_logic_vector(0 downto 0);
	signal m_p2_data_in, m_p2_data_out :
		std_logic_vector((DATA_WIDTH-1) downto 0);
	signal m_p2_addr : std_logic_vector((ADDR_WIDTH-1) downto 0);
	signal m_p2_clk, m_p2_en, m_p2_ssr, m_p2_we : std_logic;

begin

	m_p1_en <= '1';
	m_p2_en <= '1';

	m_p1_ssr <= reset;
	m_p2_ssr <= reset;

	m_p1_addr <= p1_addr;
	m_p2_addr <= p2_addr;

	p1_data_out <= m_p1_data_out;
	p2_data_out <= m_p2_data_out;

	m_p1_data_in <= p1_data_in;
	m_p2_data_in <= p2_data_in;

	m_p1_clk <= clk;
	m_p2_clk <= clk;

	m_p1_we <= p1_strobe;
	m_p2_we <= p2_strobe;

	-- RAMB16_S9_S9: Virtex-II/II-Pro, Spartan-3/3E 2k x 8 + 1 Parity bit Dual-Port RAM
	-- Xilinx HDL Language Template, version 9.1i

	RAMB16_S9_S9_inst : RAMB16_S9_S9
	generic map (
		INIT_A => X"000", --  Value of output RAM registers on Port A at startup
		INIT_B => X"000", --  Value of output RAM registers on Port B at startup
		SRVAL_A => X"000", --  Port A ouput value upon SSR assertion
		SRVAL_B => X"000", --  Port B ouput value upon SSR assertion
		WRITE_MODE_A => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
		WRITE_MODE_B => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
		SIM_COLLISION_CHECK => "ALL", -- "NONE", "WARNING", "GENERATE_X_ONLY", "ALL" 
		-- The following INIT_xx declarations specify the initial contents of the RAM
		-- Address 0 to 511
		INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
		-- Address 512 to 1023
		INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
		-- Address 1024 to 1535
		INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
		-- Address 1536 to 2047
		INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
		-- The next set of INITP_xx are for the parity bits
		-- Address 0 to 511
		INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
		-- Address 512 to 1023
		INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
		-- Address 1024 to 1535
		INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
		-- Address 1536 to 2047
		INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
	port map (
		DOA => m_p1_data_out,		-- Port A 8-bit Data Output
		DOB => m_p2_data_out,		-- Port B 8-bit Data Output
		DOPA => m_p1_parity_out,	 -- Port A 1-bit Parity Output
		DOPB => m_p2_parity_out,	 -- Port B 1-bit Parity Output
		ADDRA => m_p1_addr,  -- Port A 11-bit Address Input
		ADDRB => m_p2_addr,  -- Port B 11-bit Address Input
		CLKA => m_p1_clk,	 -- Port A Clock
		CLKB => m_p2_clk,	 -- Port B Clock
		DIA => m_p1_data_in,		-- Port A 8-bit Data Input
		DIB => m_p2_data_in,		-- Port B 8-bit Data Input
		DIPA => m_p1_parity_in,	 -- Port A 1-bit parity Input
		DIPB => m_p2_parity_in,	 -- Port-B 1-bit parity Input
		ENA => m_p1_en,		-- Port A RAM Enable Input
		ENB => m_p2_en,		-- PortB RAM Enable Input
		SSRA => m_p1_ssr,	 -- Port A Synchronous Set/Reset Input
		SSRB => m_p2_ssr,	 -- Port B Synchronous Set/Reset Input
		WEA => m_p1_we,		-- Port A Write Enable Input
		WEB => m_p2_we		 -- Port B Write Enable Input
	);

end arch;

